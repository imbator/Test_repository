library verilog;
use verilog.vl_types.all;
entity custom_reg_vlg_vec_tst is
end custom_reg_vlg_vec_tst;
