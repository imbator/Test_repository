library verilog;
use verilog.vl_types.all;
entity custom_trigger_vlg_vec_tst is
end custom_trigger_vlg_vec_tst;
